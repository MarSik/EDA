.MODEL irkd235 d
+IS=7.75629e-16 RS=0.46044 N=1.09796 EG=1.23653
+XTI=3.30648 BV=2200 IBV=0.05 CJO=1e-11
+VJ=0.7 M=0.5 FC=0.5 TT=1e-09
+KF=0 AF=1
* Model generated on Jun  3, 96
* Model format: SPICE3

