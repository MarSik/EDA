.MODEL 5eq100 d
+IS=8.77154e-05 RS=0.0202145 N=2 EG=0.815312
+XTI=3.9995 BV=100 IBV=0.005 CJO=1.06148e-09
+VJ=0.79108 M=0.475554 FC=0.5 TT=0
+KF=0 AF=1
* Model generated on May 28, 96
* Model format: SPICE3

