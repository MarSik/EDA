.MODEL 8eq045 d
+IS=1.8026e-05 RS=0.0138308 N=1.50131 EG=0.689509
+XTI=4 BV=45 IBV=0.005 CJO=1.98488e-09
+VJ=0.711167 M=0.477336 FC=0.5 TT=0
+KF=0 AF=1
* Model generated on May 28, 96
* Model format: SPICE3

